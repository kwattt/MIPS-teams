module Shift_left_J(
	input[25:0] entrada,
	output[25:0] salida

);
assign salida = {entrada<<2};

endmodule 