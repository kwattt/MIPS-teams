module Shift_left(
	input[31:0] sing_ext,
	output[31:0] salida

);

endmodule 