module Shift_left(
	input[31:0] entrada,
	output[31:0] salida

);
assign 

	salida = entrada<<32;

endmodule 